library IEEE; use IEEE.STD_LOGIC_1164.all; 
 
entity tristate is   
	port(a: in STD_LOGIC_VECTOR(15 downto 0);        
		 en: in STD_LOGIC;         
		 y: out STD_LOGIC_VECTOR(15 downto 0)); 

end;  

architecture synth of tristate is 
begin   
	y <= a when en = '1' else "ZZZZZZZZZZZZZZZZ"; 
end;   