library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_arith.ALL;
use IEEE.STD_LOGIC_unsigned.ALL;
use STD.TEXTIO.ALL ;

entity testbench_vua is -- no inputs or outputs
end;
architecture sim of testbench_vua is
	component vua
		port (p, g: in  STD_LOGIC_VECTOR(3 downto 0);
			  pg, gg: out  STD_LOGIC;
		      cin: in  STD_LOGIC;
		      c: out STD_LOGIC_VECTOR(3 downto 0));
	end component;
signal clk: STD_LOGIC;
signal p, g, c: STD_LOGIC_VECTOR(3 downto 0);
signal pg, gg: STD_LOGIC;
signal cin: STD_LOGIC;
signal pgexpected: STD_LOGIC;
Signal ggexpected: STD_LOGIC;
Signal cexpected: STD_LOGIC_VECTOR(3 downto 0);

constant MEMSIZE: integer := 32; --
type tvarray is array (MEMSIZE-1 downto 0) of
STD_LOGIC_VECTOR (14 downto 0);
signal testvectors: tvarray;
shared variable vectornum, errors: integer;
begin
-- instantiate device under test
dut: vua port map (p, g, pg, gg, cin, c);
-- generate clock
process begin
	clk <= '1'; wait for 15 ns;  
	clk <= '0'; wait for 5 ns;
end process;
-- at start of test, load vectors
-- and pulse reset
process is
file tv: TEXT;
variable i, j: integer;
variable L: line;
variable ch: character;
begin
	-- read file of test vectors
	i := 0;
	FILE_OPEN (tv, "./vua.tv", READ_MODE);
	while not endfile(tv) loop
		readline (tv, L);
		for j in 14 downto 0 loop
			read (L, ch);
			if (ch = '_') then read (L, ch);
			end if;
			if (ch = '0') then
			testvectors (i) (j) <= '0';
			else testvectors (i) (j) <= '1';
			end if;
		end loop;
		i := i + 1;
	end loop;
	vectornum := 0; errors := 0;
	-- reset <= '1'; wait for 27 ns; reset <= '0';
	wait;
end process;
-- apply test vectors on rising edge of clk
process (clk) begin
	if (clk'event and clk='1') then   
		cin <= testvectors (vectornum) (14); --after 1 ns;
		p <= testvectors (vectornum) (13 downto 10); --after 1 ns;
		g <= testvectors (vectornum) (9 downto 6); --after 1 ns;
		
		cexpected <= testvectors (vectornum)(5 downto 2); --after 1 ns;
		pgexpected <= testvectors (vectornum)(1); --after 1 ns;
		ggexpected <= testvectors (vectornum)(0); --after 1 ns;

	end if;
end process;
-- check results on falling edge of clk
process (clk) begin
	if (clk'event and clk = '0')then
		
			assert pg = pgexpected
			report "Vetor deu erro n. Teste: " &integer'image(vectornum)&". Esperado pgesp ="& STD_LOGIC'image(pgexpected)&"Valor Obtido: pg ="& STD_LOGIC'image(pg);
			if (pg /= pgexpected) then
				errors := errors + 1;
			end if;
			
			assert gg = ggexpected
			report "Vetor deu erro n. Teste: " &integer'image(vectornum)&". Esperado ggesp ="& STD_LOGIC'image(ggexpected)&"Valor Obtido: gg ="& STD_LOGIC'image(gg);
			if (gg /= ggexpected) then
			  errors := errors + 1;
			end if;  
			
			for k in 0 to 3 loop
			if(cexpected(k)='U')then
			else
				assert c(k)= cexpected(k)
					report "Vetor deu erro n. Teste: " &integer'image(vectornum)&". Esperado qesp ="& STD_LOGIC'image(cexpected(k))&"Valor Obtido: c("&integer'image(k)&") ="& STD_LOGIC'image(c(k));
				
				if (c(k)/= cexpected(k)) then
					errors := errors + 1;
				end if;
			end if;
		end loop;

			vectornum := vectornum + 1;
				  
	
		
		
		
		if (vectornum = MEMSIZE) then
			if (errors = 0) then
				report "Just kidding --" &
				integer'image (vectornum) &
				"tests completed successfully."
				severity failure;
			else
				report integer'image (vectornum) &
				"tests completed, errors = " &
				integer'image (errors)
				severity failure;
			end if;
		end if;
	end if;
	
end process;
end;
